package and2comp_pack is
	component and2
		port( a : in bit; b : in bit; c : out bit); 
	end component; 
end and2comp_pack;
